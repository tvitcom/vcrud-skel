// module main

// import vweb
// import markdown

// pub fn as_html(str string) vweb.RawHtml {
// 	return vweb.RawHtml(markdown.to_html(str))
// }